module lab1(LED, SW);
input [9:0] SW;
output [9:0] LED;

assign LED = SW;
endmodule
